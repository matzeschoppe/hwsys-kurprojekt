declare bus BUTTON1_IN, BUTTON2_IN, BUTTON3_IN, BUTTON4_IN, START_IN;
declare bus PLAYER1_BUTTON_LEFT_OUT, PLAYER1_BUTTON_RIGHT_OUT, 
	        PLAYER2_BUTTON_LEFT_OUT, PLAYER2_BUTTON_RIGHT_OUT, START_OUT;

declare register LOCKED;

RESET: 
LOCKED <- 0;
PLAYER1_BUTTON_LEFT_OUT = 0, PLAYER1_BUTTON_RIGHT_OUT = 0, 
PLAYER2_BUTTON_LEFT_OUT = 0, PLAYER2_BUTTON_RIGHT_OUT = 0, START_OUT = 0;


LOOP:
if LOCKED = 0 then 
    if BUTTON1_IN = 1 then
        PLAYER1_BUTTON_LEFT_OUT <- 1, LOCKED <- 1;
    else if BUTTON2_IN = 1 then
        PLAYER1_BUTTON_RIGHT_OUT <- 1, LOCKED <- 1;
    else if BUTTON3_IN = 1 then
        PLAYER2_BUTTON_LEFT_OUT <- 1, LOCKED <- 1;
    else if BUTTON4_IN = 1 then
        PLAYER2_BUTTON_RIGHT_OUT <- 1, LOCKED <- 1;
    fi;
fi;
if START_IN = 1 then 
    START_OUT <- 1;
    WAIT(10);
    goto RESET fi;
